`timescale 1ns / 1ps
module fpu_tb();
reg clk;
//reg opcode;
reg [15:0] A0,B0,A1,B1,A2,B2,A3,B3,A4,B4,A5,B5,A6,B6,A7,B7,A8,B8,A9,B9,A10,B10,A11,B11;
wire [15:0] dot_product;
initial begin
clk=0;
forever #5 clk=~clk;
end
MAC
uut1(clk,A0,B0,A1,B1,A2,B2,A3,B3,A4,B4,A5,B5,A6,B6,A7,B7,A8,B8,A9,B9,A10,B10,A11,B11,dot_product);
initial begin
A0 = 16'b0010111001100110;//2e66
A1 = 16'b0011001001100110;//3266
A2 = 16'b0011010000000000;//3400
A3 = 16'b1011010011001101;//b4cd
A4 = 16'b0011011001100110;//3666
A5 = 16'b0011100000000000;//3800
A6 = 16'b0011100001100110;//3866
A7 = 16'b0011100011001101;//38cd
A8 = 16'b1011101000000000;//ba00
A9 = 16'b0011101001100110;//3a66
A10 = 16'b0011101100000000;//3b00
A11 = 16'b0011101100110011;//3b33
B0 = 16'b0011010001010010;//3452
B1 = 16'b1011101110011010;//bb9a
B2 = 16'b0011000000000000;//3000
B3 = 16'b0011101001100110;//3a66
B4 = 16'b0011101100000000;//3b00
B5 = 16'b1011101000000000;//ba00
B6 = 16'b0011011001100110;//3666
B7 = 16'b0011100011001101;//38cd
B8 = 16'b0011000011001101;//30cd
B9 = 16'b0011010000000000;//3400
B10 = 16'b1011011001100110;//b666
B11 = 16'b0011100001100110;//3866
#20;
$finish;
end
endmodule
